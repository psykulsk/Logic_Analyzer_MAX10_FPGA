module Controller (
	uartMessage,
	clk_10MHz,
	fifoFull,
	fifoEmpty,
	capture,
	triggerMask,
	triggerBlockReset,
	fifoReset
	
	
	);